`ifndef RV32_CONSTS_SVH
`define RV32_CONSTS_SVH

package RV32Consts;
    localparam XLEN = 32;
    typedef logic[XLEN-1:0] IntReg;
endpackage


`endif